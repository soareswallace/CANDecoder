module can_decoder